../temp_calc_v1_0/TempCalc.vhd