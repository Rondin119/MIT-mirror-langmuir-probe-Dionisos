../set_voltage_v1_0/SetVolts.vhd