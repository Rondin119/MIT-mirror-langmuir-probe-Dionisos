../data_collector_v1_0/DataCollect.vhd