../vfloat_calc_v1_0/vFloat.vhd